// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_proj_example
 *
 * This is an example of a (trivially simple) user project,
 * showing how the user project can connect to the logic
 * analyzer, the wishbone bus, and the I/O pads.
 *
 * This project generates an integer count, which is output
 * on the user area GPIO pads (digital output only).  The
 * wishbone connection allows the project to be controlled
 * (start and stop) from the management SoC program.
 *
 * See the testbenches in directory "mprj_counter" for the
 * example programs that drive this user project.  The three
 * testbenches are "io_ports", "la_test1", and "la_test2".
 *
 *-------------------------------------------------------------
 */

 

module user_proj_datapath #(
    parameter BITS = 32
)(
`ifdef USE_POWER_PINS
    inout vccd1,	// User area 1 1.8V supply
    inout vssd1,	// User area 1 digital ground
`endif

    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,

    // IOs
    output [BITS-1:0] io_out,
    output [BITS-1:0] io_oeb,

    // Logic Analyzer Signals
    input  [127:0] la_data_in,
    output [127:0] la_data_out,
    input  [127:0] la_oenb
);

wire ALUSrc, AddSub, Cout, Overflow, clk, rst;
wire[4:0] RA0, RA1, WA;
wire[31:0] ALUout;
wire[15:0] Im;


assign clk = (~la_oenb[64]) ? la_data_in[64]: wb_clk_i;
assign rst = (~la_oenb[65]) ? la_data_in[65]: wb_rst_i;

assign {ALUSrc, AddSub, RA0, RA1, WA, Im} = la_data_in[32:0];

datapath1 datapath(
    .i_CLK(clk),
    .i_ALUSrc(ALUSrc),
    .i_AddSub(AddSub),
    .i_RST(rst),
    .i_RA0(RA0),
    .i_RA1(RA1),
    .i_WA(WA),
    .i_Im(Im),
    .o_Cout(Cout),
    .o_Overflow(Overflow),
    .o_ALUout(ALUout)
);

assign la_data_out = {ALUout, Cout, Overflow,  94'b0};
assign io_out = {ALUout};
assign io_oeb = {32'b0};

endmodule

`default_nettype wire
