magic
tech sky130A
magscale 1 2
timestamp 1730439483
<< obsli1 >>
rect 1104 2159 398820 497777
<< obsm1 >>
rect 934 552 398820 497808
<< metal2 >>
rect 5170 0 5226 800
rect 6182 0 6238 800
rect 7194 0 7250 800
rect 8206 0 8262 800
rect 9218 0 9274 800
rect 10230 0 10286 800
rect 11242 0 11298 800
rect 12254 0 12310 800
rect 13266 0 13322 800
rect 14278 0 14334 800
rect 15290 0 15346 800
rect 16302 0 16358 800
rect 17314 0 17370 800
rect 18326 0 18382 800
rect 19338 0 19394 800
rect 20350 0 20406 800
rect 21362 0 21418 800
rect 22374 0 22430 800
rect 23386 0 23442 800
rect 24398 0 24454 800
rect 25410 0 25466 800
rect 26422 0 26478 800
rect 27434 0 27490 800
rect 28446 0 28502 800
rect 29458 0 29514 800
rect 30470 0 30526 800
rect 31482 0 31538 800
rect 32494 0 32550 800
rect 33506 0 33562 800
rect 34518 0 34574 800
rect 35530 0 35586 800
rect 36542 0 36598 800
rect 37554 0 37610 800
rect 38566 0 38622 800
rect 39578 0 39634 800
rect 40590 0 40646 800
rect 41602 0 41658 800
rect 42614 0 42670 800
rect 43626 0 43682 800
rect 44638 0 44694 800
rect 45650 0 45706 800
rect 46662 0 46718 800
rect 47674 0 47730 800
rect 48686 0 48742 800
rect 49698 0 49754 800
rect 50710 0 50766 800
rect 51722 0 51778 800
rect 52734 0 52790 800
rect 53746 0 53802 800
rect 54758 0 54814 800
rect 55770 0 55826 800
rect 56782 0 56838 800
rect 57794 0 57850 800
rect 58806 0 58862 800
rect 59818 0 59874 800
rect 60830 0 60886 800
rect 61842 0 61898 800
rect 62854 0 62910 800
rect 63866 0 63922 800
rect 64878 0 64934 800
rect 65890 0 65946 800
rect 66902 0 66958 800
rect 67914 0 67970 800
rect 68926 0 68982 800
rect 69938 0 69994 800
rect 70950 0 71006 800
rect 71962 0 72018 800
rect 72974 0 73030 800
rect 73986 0 74042 800
rect 74998 0 75054 800
rect 76010 0 76066 800
rect 77022 0 77078 800
rect 78034 0 78090 800
rect 79046 0 79102 800
rect 80058 0 80114 800
rect 81070 0 81126 800
rect 82082 0 82138 800
rect 83094 0 83150 800
rect 84106 0 84162 800
rect 85118 0 85174 800
rect 86130 0 86186 800
rect 87142 0 87198 800
rect 88154 0 88210 800
rect 89166 0 89222 800
rect 90178 0 90234 800
rect 91190 0 91246 800
rect 92202 0 92258 800
rect 93214 0 93270 800
rect 94226 0 94282 800
rect 95238 0 95294 800
rect 96250 0 96306 800
rect 97262 0 97318 800
rect 98274 0 98330 800
rect 99286 0 99342 800
rect 100298 0 100354 800
rect 101310 0 101366 800
rect 102322 0 102378 800
rect 103334 0 103390 800
rect 104346 0 104402 800
rect 105358 0 105414 800
rect 106370 0 106426 800
rect 107382 0 107438 800
rect 108394 0 108450 800
rect 109406 0 109462 800
rect 110418 0 110474 800
rect 111430 0 111486 800
rect 112442 0 112498 800
rect 113454 0 113510 800
rect 114466 0 114522 800
rect 115478 0 115534 800
rect 116490 0 116546 800
rect 117502 0 117558 800
rect 118514 0 118570 800
rect 119526 0 119582 800
rect 120538 0 120594 800
rect 121550 0 121606 800
rect 122562 0 122618 800
rect 123574 0 123630 800
rect 124586 0 124642 800
rect 125598 0 125654 800
rect 126610 0 126666 800
rect 127622 0 127678 800
rect 128634 0 128690 800
rect 129646 0 129702 800
rect 130658 0 130714 800
rect 131670 0 131726 800
rect 132682 0 132738 800
rect 133694 0 133750 800
rect 134706 0 134762 800
rect 135718 0 135774 800
rect 136730 0 136786 800
rect 137742 0 137798 800
rect 138754 0 138810 800
rect 139766 0 139822 800
rect 140778 0 140834 800
rect 141790 0 141846 800
rect 142802 0 142858 800
rect 143814 0 143870 800
rect 144826 0 144882 800
rect 145838 0 145894 800
rect 146850 0 146906 800
rect 147862 0 147918 800
rect 148874 0 148930 800
rect 149886 0 149942 800
rect 150898 0 150954 800
rect 151910 0 151966 800
rect 152922 0 152978 800
rect 153934 0 153990 800
rect 154946 0 155002 800
rect 155958 0 156014 800
rect 156970 0 157026 800
rect 157982 0 158038 800
rect 158994 0 159050 800
rect 160006 0 160062 800
rect 161018 0 161074 800
rect 162030 0 162086 800
rect 163042 0 163098 800
rect 164054 0 164110 800
rect 165066 0 165122 800
rect 166078 0 166134 800
rect 167090 0 167146 800
rect 168102 0 168158 800
rect 169114 0 169170 800
rect 170126 0 170182 800
rect 171138 0 171194 800
rect 172150 0 172206 800
rect 173162 0 173218 800
rect 174174 0 174230 800
rect 175186 0 175242 800
rect 176198 0 176254 800
rect 177210 0 177266 800
rect 178222 0 178278 800
rect 179234 0 179290 800
rect 180246 0 180302 800
rect 181258 0 181314 800
rect 182270 0 182326 800
rect 183282 0 183338 800
rect 184294 0 184350 800
rect 185306 0 185362 800
rect 186318 0 186374 800
rect 187330 0 187386 800
rect 188342 0 188398 800
rect 189354 0 189410 800
rect 190366 0 190422 800
rect 191378 0 191434 800
rect 192390 0 192446 800
rect 193402 0 193458 800
rect 194414 0 194470 800
rect 195426 0 195482 800
rect 196438 0 196494 800
rect 197450 0 197506 800
rect 198462 0 198518 800
rect 199474 0 199530 800
rect 200486 0 200542 800
rect 201498 0 201554 800
rect 202510 0 202566 800
rect 203522 0 203578 800
rect 204534 0 204590 800
rect 205546 0 205602 800
rect 206558 0 206614 800
rect 207570 0 207626 800
rect 208582 0 208638 800
rect 209594 0 209650 800
rect 210606 0 210662 800
rect 211618 0 211674 800
rect 212630 0 212686 800
rect 213642 0 213698 800
rect 214654 0 214710 800
rect 215666 0 215722 800
rect 216678 0 216734 800
rect 217690 0 217746 800
rect 218702 0 218758 800
rect 219714 0 219770 800
rect 220726 0 220782 800
rect 221738 0 221794 800
rect 222750 0 222806 800
rect 223762 0 223818 800
rect 224774 0 224830 800
rect 225786 0 225842 800
rect 226798 0 226854 800
rect 227810 0 227866 800
rect 228822 0 228878 800
rect 229834 0 229890 800
rect 230846 0 230902 800
rect 231858 0 231914 800
rect 232870 0 232926 800
rect 233882 0 233938 800
rect 234894 0 234950 800
rect 235906 0 235962 800
rect 236918 0 236974 800
rect 237930 0 237986 800
rect 238942 0 238998 800
rect 239954 0 240010 800
rect 240966 0 241022 800
rect 241978 0 242034 800
rect 242990 0 243046 800
rect 244002 0 244058 800
rect 245014 0 245070 800
rect 246026 0 246082 800
rect 247038 0 247094 800
rect 248050 0 248106 800
rect 249062 0 249118 800
rect 250074 0 250130 800
rect 251086 0 251142 800
rect 252098 0 252154 800
rect 253110 0 253166 800
rect 254122 0 254178 800
rect 255134 0 255190 800
rect 256146 0 256202 800
rect 257158 0 257214 800
rect 258170 0 258226 800
rect 259182 0 259238 800
rect 260194 0 260250 800
rect 261206 0 261262 800
rect 262218 0 262274 800
rect 263230 0 263286 800
rect 264242 0 264298 800
rect 265254 0 265310 800
rect 266266 0 266322 800
rect 267278 0 267334 800
rect 268290 0 268346 800
rect 269302 0 269358 800
rect 270314 0 270370 800
rect 271326 0 271382 800
rect 272338 0 272394 800
rect 273350 0 273406 800
rect 274362 0 274418 800
rect 275374 0 275430 800
rect 276386 0 276442 800
rect 277398 0 277454 800
rect 278410 0 278466 800
rect 279422 0 279478 800
rect 280434 0 280490 800
rect 281446 0 281502 800
rect 282458 0 282514 800
rect 283470 0 283526 800
rect 284482 0 284538 800
rect 285494 0 285550 800
rect 286506 0 286562 800
rect 287518 0 287574 800
rect 288530 0 288586 800
rect 289542 0 289598 800
rect 290554 0 290610 800
rect 291566 0 291622 800
rect 292578 0 292634 800
rect 293590 0 293646 800
rect 294602 0 294658 800
rect 295614 0 295670 800
rect 296626 0 296682 800
rect 297638 0 297694 800
rect 298650 0 298706 800
rect 299662 0 299718 800
rect 300674 0 300730 800
rect 301686 0 301742 800
rect 302698 0 302754 800
rect 303710 0 303766 800
rect 304722 0 304778 800
rect 305734 0 305790 800
rect 306746 0 306802 800
rect 307758 0 307814 800
rect 308770 0 308826 800
rect 309782 0 309838 800
rect 310794 0 310850 800
rect 311806 0 311862 800
rect 312818 0 312874 800
rect 313830 0 313886 800
rect 314842 0 314898 800
rect 315854 0 315910 800
rect 316866 0 316922 800
rect 317878 0 317934 800
rect 318890 0 318946 800
rect 319902 0 319958 800
rect 320914 0 320970 800
rect 321926 0 321982 800
rect 322938 0 322994 800
rect 323950 0 324006 800
rect 324962 0 325018 800
rect 325974 0 326030 800
rect 326986 0 327042 800
rect 327998 0 328054 800
rect 329010 0 329066 800
rect 330022 0 330078 800
rect 331034 0 331090 800
rect 332046 0 332102 800
rect 333058 0 333114 800
rect 334070 0 334126 800
rect 335082 0 335138 800
rect 336094 0 336150 800
rect 337106 0 337162 800
rect 338118 0 338174 800
rect 339130 0 339186 800
rect 340142 0 340198 800
rect 341154 0 341210 800
rect 342166 0 342222 800
rect 343178 0 343234 800
rect 344190 0 344246 800
rect 345202 0 345258 800
rect 346214 0 346270 800
rect 347226 0 347282 800
rect 348238 0 348294 800
rect 349250 0 349306 800
rect 350262 0 350318 800
rect 351274 0 351330 800
rect 352286 0 352342 800
rect 353298 0 353354 800
rect 354310 0 354366 800
rect 355322 0 355378 800
rect 356334 0 356390 800
rect 357346 0 357402 800
rect 358358 0 358414 800
rect 359370 0 359426 800
rect 360382 0 360438 800
rect 361394 0 361450 800
rect 362406 0 362462 800
rect 363418 0 363474 800
rect 364430 0 364486 800
rect 365442 0 365498 800
rect 366454 0 366510 800
rect 367466 0 367522 800
rect 368478 0 368534 800
rect 369490 0 369546 800
rect 370502 0 370558 800
rect 371514 0 371570 800
rect 372526 0 372582 800
rect 373538 0 373594 800
rect 374550 0 374606 800
rect 375562 0 375618 800
rect 376574 0 376630 800
rect 377586 0 377642 800
rect 378598 0 378654 800
rect 379610 0 379666 800
rect 380622 0 380678 800
rect 381634 0 381690 800
rect 382646 0 382702 800
rect 383658 0 383714 800
rect 384670 0 384726 800
rect 385682 0 385738 800
rect 386694 0 386750 800
rect 387706 0 387762 800
rect 388718 0 388774 800
rect 389730 0 389786 800
rect 390742 0 390798 800
rect 391754 0 391810 800
rect 392766 0 392822 800
rect 393778 0 393834 800
rect 394790 0 394846 800
<< obsm2 >>
rect 938 856 398526 497797
rect 938 546 5114 856
rect 5282 546 6126 856
rect 6294 546 7138 856
rect 7306 546 8150 856
rect 8318 546 9162 856
rect 9330 546 10174 856
rect 10342 546 11186 856
rect 11354 546 12198 856
rect 12366 546 13210 856
rect 13378 546 14222 856
rect 14390 546 15234 856
rect 15402 546 16246 856
rect 16414 546 17258 856
rect 17426 546 18270 856
rect 18438 546 19282 856
rect 19450 546 20294 856
rect 20462 546 21306 856
rect 21474 546 22318 856
rect 22486 546 23330 856
rect 23498 546 24342 856
rect 24510 546 25354 856
rect 25522 546 26366 856
rect 26534 546 27378 856
rect 27546 546 28390 856
rect 28558 546 29402 856
rect 29570 546 30414 856
rect 30582 546 31426 856
rect 31594 546 32438 856
rect 32606 546 33450 856
rect 33618 546 34462 856
rect 34630 546 35474 856
rect 35642 546 36486 856
rect 36654 546 37498 856
rect 37666 546 38510 856
rect 38678 546 39522 856
rect 39690 546 40534 856
rect 40702 546 41546 856
rect 41714 546 42558 856
rect 42726 546 43570 856
rect 43738 546 44582 856
rect 44750 546 45594 856
rect 45762 546 46606 856
rect 46774 546 47618 856
rect 47786 546 48630 856
rect 48798 546 49642 856
rect 49810 546 50654 856
rect 50822 546 51666 856
rect 51834 546 52678 856
rect 52846 546 53690 856
rect 53858 546 54702 856
rect 54870 546 55714 856
rect 55882 546 56726 856
rect 56894 546 57738 856
rect 57906 546 58750 856
rect 58918 546 59762 856
rect 59930 546 60774 856
rect 60942 546 61786 856
rect 61954 546 62798 856
rect 62966 546 63810 856
rect 63978 546 64822 856
rect 64990 546 65834 856
rect 66002 546 66846 856
rect 67014 546 67858 856
rect 68026 546 68870 856
rect 69038 546 69882 856
rect 70050 546 70894 856
rect 71062 546 71906 856
rect 72074 546 72918 856
rect 73086 546 73930 856
rect 74098 546 74942 856
rect 75110 546 75954 856
rect 76122 546 76966 856
rect 77134 546 77978 856
rect 78146 546 78990 856
rect 79158 546 80002 856
rect 80170 546 81014 856
rect 81182 546 82026 856
rect 82194 546 83038 856
rect 83206 546 84050 856
rect 84218 546 85062 856
rect 85230 546 86074 856
rect 86242 546 87086 856
rect 87254 546 88098 856
rect 88266 546 89110 856
rect 89278 546 90122 856
rect 90290 546 91134 856
rect 91302 546 92146 856
rect 92314 546 93158 856
rect 93326 546 94170 856
rect 94338 546 95182 856
rect 95350 546 96194 856
rect 96362 546 97206 856
rect 97374 546 98218 856
rect 98386 546 99230 856
rect 99398 546 100242 856
rect 100410 546 101254 856
rect 101422 546 102266 856
rect 102434 546 103278 856
rect 103446 546 104290 856
rect 104458 546 105302 856
rect 105470 546 106314 856
rect 106482 546 107326 856
rect 107494 546 108338 856
rect 108506 546 109350 856
rect 109518 546 110362 856
rect 110530 546 111374 856
rect 111542 546 112386 856
rect 112554 546 113398 856
rect 113566 546 114410 856
rect 114578 546 115422 856
rect 115590 546 116434 856
rect 116602 546 117446 856
rect 117614 546 118458 856
rect 118626 546 119470 856
rect 119638 546 120482 856
rect 120650 546 121494 856
rect 121662 546 122506 856
rect 122674 546 123518 856
rect 123686 546 124530 856
rect 124698 546 125542 856
rect 125710 546 126554 856
rect 126722 546 127566 856
rect 127734 546 128578 856
rect 128746 546 129590 856
rect 129758 546 130602 856
rect 130770 546 131614 856
rect 131782 546 132626 856
rect 132794 546 133638 856
rect 133806 546 134650 856
rect 134818 546 135662 856
rect 135830 546 136674 856
rect 136842 546 137686 856
rect 137854 546 138698 856
rect 138866 546 139710 856
rect 139878 546 140722 856
rect 140890 546 141734 856
rect 141902 546 142746 856
rect 142914 546 143758 856
rect 143926 546 144770 856
rect 144938 546 145782 856
rect 145950 546 146794 856
rect 146962 546 147806 856
rect 147974 546 148818 856
rect 148986 546 149830 856
rect 149998 546 150842 856
rect 151010 546 151854 856
rect 152022 546 152866 856
rect 153034 546 153878 856
rect 154046 546 154890 856
rect 155058 546 155902 856
rect 156070 546 156914 856
rect 157082 546 157926 856
rect 158094 546 158938 856
rect 159106 546 159950 856
rect 160118 546 160962 856
rect 161130 546 161974 856
rect 162142 546 162986 856
rect 163154 546 163998 856
rect 164166 546 165010 856
rect 165178 546 166022 856
rect 166190 546 167034 856
rect 167202 546 168046 856
rect 168214 546 169058 856
rect 169226 546 170070 856
rect 170238 546 171082 856
rect 171250 546 172094 856
rect 172262 546 173106 856
rect 173274 546 174118 856
rect 174286 546 175130 856
rect 175298 546 176142 856
rect 176310 546 177154 856
rect 177322 546 178166 856
rect 178334 546 179178 856
rect 179346 546 180190 856
rect 180358 546 181202 856
rect 181370 546 182214 856
rect 182382 546 183226 856
rect 183394 546 184238 856
rect 184406 546 185250 856
rect 185418 546 186262 856
rect 186430 546 187274 856
rect 187442 546 188286 856
rect 188454 546 189298 856
rect 189466 546 190310 856
rect 190478 546 191322 856
rect 191490 546 192334 856
rect 192502 546 193346 856
rect 193514 546 194358 856
rect 194526 546 195370 856
rect 195538 546 196382 856
rect 196550 546 197394 856
rect 197562 546 198406 856
rect 198574 546 199418 856
rect 199586 546 200430 856
rect 200598 546 201442 856
rect 201610 546 202454 856
rect 202622 546 203466 856
rect 203634 546 204478 856
rect 204646 546 205490 856
rect 205658 546 206502 856
rect 206670 546 207514 856
rect 207682 546 208526 856
rect 208694 546 209538 856
rect 209706 546 210550 856
rect 210718 546 211562 856
rect 211730 546 212574 856
rect 212742 546 213586 856
rect 213754 546 214598 856
rect 214766 546 215610 856
rect 215778 546 216622 856
rect 216790 546 217634 856
rect 217802 546 218646 856
rect 218814 546 219658 856
rect 219826 546 220670 856
rect 220838 546 221682 856
rect 221850 546 222694 856
rect 222862 546 223706 856
rect 223874 546 224718 856
rect 224886 546 225730 856
rect 225898 546 226742 856
rect 226910 546 227754 856
rect 227922 546 228766 856
rect 228934 546 229778 856
rect 229946 546 230790 856
rect 230958 546 231802 856
rect 231970 546 232814 856
rect 232982 546 233826 856
rect 233994 546 234838 856
rect 235006 546 235850 856
rect 236018 546 236862 856
rect 237030 546 237874 856
rect 238042 546 238886 856
rect 239054 546 239898 856
rect 240066 546 240910 856
rect 241078 546 241922 856
rect 242090 546 242934 856
rect 243102 546 243946 856
rect 244114 546 244958 856
rect 245126 546 245970 856
rect 246138 546 246982 856
rect 247150 546 247994 856
rect 248162 546 249006 856
rect 249174 546 250018 856
rect 250186 546 251030 856
rect 251198 546 252042 856
rect 252210 546 253054 856
rect 253222 546 254066 856
rect 254234 546 255078 856
rect 255246 546 256090 856
rect 256258 546 257102 856
rect 257270 546 258114 856
rect 258282 546 259126 856
rect 259294 546 260138 856
rect 260306 546 261150 856
rect 261318 546 262162 856
rect 262330 546 263174 856
rect 263342 546 264186 856
rect 264354 546 265198 856
rect 265366 546 266210 856
rect 266378 546 267222 856
rect 267390 546 268234 856
rect 268402 546 269246 856
rect 269414 546 270258 856
rect 270426 546 271270 856
rect 271438 546 272282 856
rect 272450 546 273294 856
rect 273462 546 274306 856
rect 274474 546 275318 856
rect 275486 546 276330 856
rect 276498 546 277342 856
rect 277510 546 278354 856
rect 278522 546 279366 856
rect 279534 546 280378 856
rect 280546 546 281390 856
rect 281558 546 282402 856
rect 282570 546 283414 856
rect 283582 546 284426 856
rect 284594 546 285438 856
rect 285606 546 286450 856
rect 286618 546 287462 856
rect 287630 546 288474 856
rect 288642 546 289486 856
rect 289654 546 290498 856
rect 290666 546 291510 856
rect 291678 546 292522 856
rect 292690 546 293534 856
rect 293702 546 294546 856
rect 294714 546 295558 856
rect 295726 546 296570 856
rect 296738 546 297582 856
rect 297750 546 298594 856
rect 298762 546 299606 856
rect 299774 546 300618 856
rect 300786 546 301630 856
rect 301798 546 302642 856
rect 302810 546 303654 856
rect 303822 546 304666 856
rect 304834 546 305678 856
rect 305846 546 306690 856
rect 306858 546 307702 856
rect 307870 546 308714 856
rect 308882 546 309726 856
rect 309894 546 310738 856
rect 310906 546 311750 856
rect 311918 546 312762 856
rect 312930 546 313774 856
rect 313942 546 314786 856
rect 314954 546 315798 856
rect 315966 546 316810 856
rect 316978 546 317822 856
rect 317990 546 318834 856
rect 319002 546 319846 856
rect 320014 546 320858 856
rect 321026 546 321870 856
rect 322038 546 322882 856
rect 323050 546 323894 856
rect 324062 546 324906 856
rect 325074 546 325918 856
rect 326086 546 326930 856
rect 327098 546 327942 856
rect 328110 546 328954 856
rect 329122 546 329966 856
rect 330134 546 330978 856
rect 331146 546 331990 856
rect 332158 546 333002 856
rect 333170 546 334014 856
rect 334182 546 335026 856
rect 335194 546 336038 856
rect 336206 546 337050 856
rect 337218 546 338062 856
rect 338230 546 339074 856
rect 339242 546 340086 856
rect 340254 546 341098 856
rect 341266 546 342110 856
rect 342278 546 343122 856
rect 343290 546 344134 856
rect 344302 546 345146 856
rect 345314 546 346158 856
rect 346326 546 347170 856
rect 347338 546 348182 856
rect 348350 546 349194 856
rect 349362 546 350206 856
rect 350374 546 351218 856
rect 351386 546 352230 856
rect 352398 546 353242 856
rect 353410 546 354254 856
rect 354422 546 355266 856
rect 355434 546 356278 856
rect 356446 546 357290 856
rect 357458 546 358302 856
rect 358470 546 359314 856
rect 359482 546 360326 856
rect 360494 546 361338 856
rect 361506 546 362350 856
rect 362518 546 363362 856
rect 363530 546 364374 856
rect 364542 546 365386 856
rect 365554 546 366398 856
rect 366566 546 367410 856
rect 367578 546 368422 856
rect 368590 546 369434 856
rect 369602 546 370446 856
rect 370614 546 371458 856
rect 371626 546 372470 856
rect 372638 546 373482 856
rect 373650 546 374494 856
rect 374662 546 375506 856
rect 375674 546 376518 856
rect 376686 546 377530 856
rect 377698 546 378542 856
rect 378710 546 379554 856
rect 379722 546 380566 856
rect 380734 546 381578 856
rect 381746 546 382590 856
rect 382758 546 383602 856
rect 383770 546 384614 856
rect 384782 546 385626 856
rect 385794 546 386638 856
rect 386806 546 387650 856
rect 387818 546 388662 856
rect 388830 546 389674 856
rect 389842 546 390686 856
rect 390854 546 391698 856
rect 391866 546 392710 856
rect 392878 546 393722 856
rect 393890 546 394734 856
rect 394902 546 398526 856
<< metal3 >>
rect 0 490152 800 490272
rect 399200 490152 400000 490272
rect 0 474648 800 474768
rect 399200 474648 400000 474768
rect 0 459144 800 459264
rect 399200 459144 400000 459264
rect 0 443640 800 443760
rect 399200 443640 400000 443760
rect 0 428136 800 428256
rect 399200 428136 400000 428256
rect 0 412632 800 412752
rect 399200 412632 400000 412752
rect 0 397128 800 397248
rect 399200 397128 400000 397248
rect 0 381624 800 381744
rect 399200 381624 400000 381744
rect 0 366120 800 366240
rect 399200 366120 400000 366240
rect 0 350616 800 350736
rect 399200 350616 400000 350736
rect 0 335112 800 335232
rect 399200 335112 400000 335232
rect 0 319608 800 319728
rect 399200 319608 400000 319728
rect 0 304104 800 304224
rect 399200 304104 400000 304224
rect 0 288600 800 288720
rect 399200 288600 400000 288720
rect 0 273096 800 273216
rect 399200 273096 400000 273216
rect 0 257592 800 257712
rect 399200 257592 400000 257712
rect 0 242088 800 242208
rect 399200 242088 400000 242208
rect 0 226584 800 226704
rect 399200 226584 400000 226704
rect 0 211080 800 211200
rect 399200 211080 400000 211200
rect 0 195576 800 195696
rect 399200 195576 400000 195696
rect 0 180072 800 180192
rect 399200 180072 400000 180192
rect 0 164568 800 164688
rect 399200 164568 400000 164688
rect 0 149064 800 149184
rect 399200 149064 400000 149184
rect 0 133560 800 133680
rect 399200 133560 400000 133680
rect 0 118056 800 118176
rect 399200 118056 400000 118176
rect 0 102552 800 102672
rect 399200 102552 400000 102672
rect 0 87048 800 87168
rect 399200 87048 400000 87168
rect 0 71544 800 71664
rect 399200 71544 400000 71664
rect 0 56040 800 56160
rect 399200 56040 400000 56160
rect 0 40536 800 40656
rect 399200 40536 400000 40656
rect 0 25032 800 25152
rect 399200 25032 400000 25152
rect 0 9528 800 9648
rect 399200 9528 400000 9648
<< obsm3 >>
rect 798 490352 399200 497793
rect 880 490072 399120 490352
rect 798 474848 399200 490072
rect 880 474568 399120 474848
rect 798 459344 399200 474568
rect 880 459064 399120 459344
rect 798 443840 399200 459064
rect 880 443560 399120 443840
rect 798 428336 399200 443560
rect 880 428056 399120 428336
rect 798 412832 399200 428056
rect 880 412552 399120 412832
rect 798 397328 399200 412552
rect 880 397048 399120 397328
rect 798 381824 399200 397048
rect 880 381544 399120 381824
rect 798 366320 399200 381544
rect 880 366040 399120 366320
rect 798 350816 399200 366040
rect 880 350536 399120 350816
rect 798 335312 399200 350536
rect 880 335032 399120 335312
rect 798 319808 399200 335032
rect 880 319528 399120 319808
rect 798 304304 399200 319528
rect 880 304024 399120 304304
rect 798 288800 399200 304024
rect 880 288520 399120 288800
rect 798 273296 399200 288520
rect 880 273016 399120 273296
rect 798 257792 399200 273016
rect 880 257512 399120 257792
rect 798 242288 399200 257512
rect 880 242008 399120 242288
rect 798 226784 399200 242008
rect 880 226504 399120 226784
rect 798 211280 399200 226504
rect 880 211000 399120 211280
rect 798 195776 399200 211000
rect 880 195496 399120 195776
rect 798 180272 399200 195496
rect 880 179992 399120 180272
rect 798 164768 399200 179992
rect 880 164488 399120 164768
rect 798 149264 399200 164488
rect 880 148984 399120 149264
rect 798 133760 399200 148984
rect 880 133480 399120 133760
rect 798 118256 399200 133480
rect 880 117976 399120 118256
rect 798 102752 399200 117976
rect 880 102472 399120 102752
rect 798 87248 399200 102472
rect 880 86968 399120 87248
rect 798 71744 399200 86968
rect 880 71464 399120 71744
rect 798 56240 399200 71464
rect 880 55960 399120 56240
rect 798 40736 399200 55960
rect 880 40456 399120 40736
rect 798 25232 399200 40456
rect 880 24952 399120 25232
rect 798 9728 399200 24952
rect 880 9448 399120 9728
rect 798 444 399200 9448
<< metal4 >>
rect 4208 2128 4528 497808
rect 19568 2128 19888 497808
rect 34928 2128 35248 497808
rect 50288 2128 50608 497808
rect 65648 2128 65968 497808
rect 81008 2128 81328 497808
rect 96368 2128 96688 497808
rect 111728 2128 112048 497808
rect 127088 2128 127408 497808
rect 142448 2128 142768 497808
rect 157808 2128 158128 497808
rect 173168 2128 173488 497808
rect 188528 2128 188848 497808
rect 203888 2128 204208 497808
rect 219248 2128 219568 497808
rect 234608 2128 234928 497808
rect 249968 2128 250288 497808
rect 265328 2128 265648 497808
rect 280688 2128 281008 497808
rect 296048 2128 296368 497808
rect 311408 2128 311728 497808
rect 326768 2128 327088 497808
rect 342128 2128 342448 497808
rect 357488 2128 357808 497808
rect 372848 2128 373168 497808
rect 388208 2128 388528 497808
<< obsm4 >>
rect 64459 2048 65568 320109
rect 66048 2048 80928 320109
rect 81408 2048 96288 320109
rect 96768 2048 111648 320109
rect 112128 2048 113285 320109
rect 64459 443 113285 2048
<< labels >>
rlabel metal3 s 399200 25032 400000 25152 6 io_oeb[0]
port 1 nsew signal output
rlabel metal3 s 399200 335112 400000 335232 6 io_oeb[10]
port 2 nsew signal output
rlabel metal3 s 399200 366120 400000 366240 6 io_oeb[11]
port 3 nsew signal output
rlabel metal3 s 399200 397128 400000 397248 6 io_oeb[12]
port 4 nsew signal output
rlabel metal3 s 399200 428136 400000 428256 6 io_oeb[13]
port 5 nsew signal output
rlabel metal3 s 399200 459144 400000 459264 6 io_oeb[14]
port 6 nsew signal output
rlabel metal3 s 399200 490152 400000 490272 6 io_oeb[15]
port 7 nsew signal output
rlabel metal3 s 0 474648 800 474768 6 io_oeb[16]
port 8 nsew signal output
rlabel metal3 s 0 443640 800 443760 6 io_oeb[17]
port 9 nsew signal output
rlabel metal3 s 0 412632 800 412752 6 io_oeb[18]
port 10 nsew signal output
rlabel metal3 s 0 381624 800 381744 6 io_oeb[19]
port 11 nsew signal output
rlabel metal3 s 399200 56040 400000 56160 6 io_oeb[1]
port 12 nsew signal output
rlabel metal3 s 0 350616 800 350736 6 io_oeb[20]
port 13 nsew signal output
rlabel metal3 s 0 319608 800 319728 6 io_oeb[21]
port 14 nsew signal output
rlabel metal3 s 0 288600 800 288720 6 io_oeb[22]
port 15 nsew signal output
rlabel metal3 s 0 257592 800 257712 6 io_oeb[23]
port 16 nsew signal output
rlabel metal3 s 0 226584 800 226704 6 io_oeb[24]
port 17 nsew signal output
rlabel metal3 s 0 195576 800 195696 6 io_oeb[25]
port 18 nsew signal output
rlabel metal3 s 0 164568 800 164688 6 io_oeb[26]
port 19 nsew signal output
rlabel metal3 s 0 133560 800 133680 6 io_oeb[27]
port 20 nsew signal output
rlabel metal3 s 0 102552 800 102672 6 io_oeb[28]
port 21 nsew signal output
rlabel metal3 s 0 71544 800 71664 6 io_oeb[29]
port 22 nsew signal output
rlabel metal3 s 399200 87048 400000 87168 6 io_oeb[2]
port 23 nsew signal output
rlabel metal3 s 0 40536 800 40656 6 io_oeb[30]
port 24 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 io_oeb[31]
port 25 nsew signal output
rlabel metal3 s 399200 118056 400000 118176 6 io_oeb[3]
port 26 nsew signal output
rlabel metal3 s 399200 149064 400000 149184 6 io_oeb[4]
port 27 nsew signal output
rlabel metal3 s 399200 180072 400000 180192 6 io_oeb[5]
port 28 nsew signal output
rlabel metal3 s 399200 211080 400000 211200 6 io_oeb[6]
port 29 nsew signal output
rlabel metal3 s 399200 242088 400000 242208 6 io_oeb[7]
port 30 nsew signal output
rlabel metal3 s 399200 273096 400000 273216 6 io_oeb[8]
port 31 nsew signal output
rlabel metal3 s 399200 304104 400000 304224 6 io_oeb[9]
port 32 nsew signal output
rlabel metal3 s 399200 9528 400000 9648 6 io_out[0]
port 33 nsew signal output
rlabel metal3 s 399200 319608 400000 319728 6 io_out[10]
port 34 nsew signal output
rlabel metal3 s 399200 350616 400000 350736 6 io_out[11]
port 35 nsew signal output
rlabel metal3 s 399200 381624 400000 381744 6 io_out[12]
port 36 nsew signal output
rlabel metal3 s 399200 412632 400000 412752 6 io_out[13]
port 37 nsew signal output
rlabel metal3 s 399200 443640 400000 443760 6 io_out[14]
port 38 nsew signal output
rlabel metal3 s 399200 474648 400000 474768 6 io_out[15]
port 39 nsew signal output
rlabel metal3 s 0 490152 800 490272 6 io_out[16]
port 40 nsew signal output
rlabel metal3 s 0 459144 800 459264 6 io_out[17]
port 41 nsew signal output
rlabel metal3 s 0 428136 800 428256 6 io_out[18]
port 42 nsew signal output
rlabel metal3 s 0 397128 800 397248 6 io_out[19]
port 43 nsew signal output
rlabel metal3 s 399200 40536 400000 40656 6 io_out[1]
port 44 nsew signal output
rlabel metal3 s 0 366120 800 366240 6 io_out[20]
port 45 nsew signal output
rlabel metal3 s 0 335112 800 335232 6 io_out[21]
port 46 nsew signal output
rlabel metal3 s 0 304104 800 304224 6 io_out[22]
port 47 nsew signal output
rlabel metal3 s 0 273096 800 273216 6 io_out[23]
port 48 nsew signal output
rlabel metal3 s 0 242088 800 242208 6 io_out[24]
port 49 nsew signal output
rlabel metal3 s 0 211080 800 211200 6 io_out[25]
port 50 nsew signal output
rlabel metal3 s 0 180072 800 180192 6 io_out[26]
port 51 nsew signal output
rlabel metal3 s 0 149064 800 149184 6 io_out[27]
port 52 nsew signal output
rlabel metal3 s 0 118056 800 118176 6 io_out[28]
port 53 nsew signal output
rlabel metal3 s 0 87048 800 87168 6 io_out[29]
port 54 nsew signal output
rlabel metal3 s 399200 71544 400000 71664 6 io_out[2]
port 55 nsew signal output
rlabel metal3 s 0 56040 800 56160 6 io_out[30]
port 56 nsew signal output
rlabel metal3 s 0 25032 800 25152 6 io_out[31]
port 57 nsew signal output
rlabel metal3 s 399200 102552 400000 102672 6 io_out[3]
port 58 nsew signal output
rlabel metal3 s 399200 133560 400000 133680 6 io_out[4]
port 59 nsew signal output
rlabel metal3 s 399200 164568 400000 164688 6 io_out[5]
port 60 nsew signal output
rlabel metal3 s 399200 195576 400000 195696 6 io_out[6]
port 61 nsew signal output
rlabel metal3 s 399200 226584 400000 226704 6 io_out[7]
port 62 nsew signal output
rlabel metal3 s 399200 257592 400000 257712 6 io_out[8]
port 63 nsew signal output
rlabel metal3 s 399200 288600 400000 288720 6 io_out[9]
port 64 nsew signal output
rlabel metal2 s 7194 0 7250 800 6 la_data_in[0]
port 65 nsew signal input
rlabel metal2 s 310794 0 310850 800 6 la_data_in[100]
port 66 nsew signal input
rlabel metal2 s 313830 0 313886 800 6 la_data_in[101]
port 67 nsew signal input
rlabel metal2 s 316866 0 316922 800 6 la_data_in[102]
port 68 nsew signal input
rlabel metal2 s 319902 0 319958 800 6 la_data_in[103]
port 69 nsew signal input
rlabel metal2 s 322938 0 322994 800 6 la_data_in[104]
port 70 nsew signal input
rlabel metal2 s 325974 0 326030 800 6 la_data_in[105]
port 71 nsew signal input
rlabel metal2 s 329010 0 329066 800 6 la_data_in[106]
port 72 nsew signal input
rlabel metal2 s 332046 0 332102 800 6 la_data_in[107]
port 73 nsew signal input
rlabel metal2 s 335082 0 335138 800 6 la_data_in[108]
port 74 nsew signal input
rlabel metal2 s 338118 0 338174 800 6 la_data_in[109]
port 75 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 la_data_in[10]
port 76 nsew signal input
rlabel metal2 s 341154 0 341210 800 6 la_data_in[110]
port 77 nsew signal input
rlabel metal2 s 344190 0 344246 800 6 la_data_in[111]
port 78 nsew signal input
rlabel metal2 s 347226 0 347282 800 6 la_data_in[112]
port 79 nsew signal input
rlabel metal2 s 350262 0 350318 800 6 la_data_in[113]
port 80 nsew signal input
rlabel metal2 s 353298 0 353354 800 6 la_data_in[114]
port 81 nsew signal input
rlabel metal2 s 356334 0 356390 800 6 la_data_in[115]
port 82 nsew signal input
rlabel metal2 s 359370 0 359426 800 6 la_data_in[116]
port 83 nsew signal input
rlabel metal2 s 362406 0 362462 800 6 la_data_in[117]
port 84 nsew signal input
rlabel metal2 s 365442 0 365498 800 6 la_data_in[118]
port 85 nsew signal input
rlabel metal2 s 368478 0 368534 800 6 la_data_in[119]
port 86 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 la_data_in[11]
port 87 nsew signal input
rlabel metal2 s 371514 0 371570 800 6 la_data_in[120]
port 88 nsew signal input
rlabel metal2 s 374550 0 374606 800 6 la_data_in[121]
port 89 nsew signal input
rlabel metal2 s 377586 0 377642 800 6 la_data_in[122]
port 90 nsew signal input
rlabel metal2 s 380622 0 380678 800 6 la_data_in[123]
port 91 nsew signal input
rlabel metal2 s 383658 0 383714 800 6 la_data_in[124]
port 92 nsew signal input
rlabel metal2 s 386694 0 386750 800 6 la_data_in[125]
port 93 nsew signal input
rlabel metal2 s 389730 0 389786 800 6 la_data_in[126]
port 94 nsew signal input
rlabel metal2 s 392766 0 392822 800 6 la_data_in[127]
port 95 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 la_data_in[12]
port 96 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_data_in[13]
port 97 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_data_in[14]
port 98 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 la_data_in[15]
port 99 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 la_data_in[16]
port 100 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_data_in[17]
port 101 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 la_data_in[18]
port 102 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 la_data_in[19]
port 103 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 la_data_in[1]
port 104 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 la_data_in[20]
port 105 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_data_in[21]
port 106 nsew signal input
rlabel metal2 s 73986 0 74042 800 6 la_data_in[22]
port 107 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 la_data_in[23]
port 108 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 la_data_in[24]
port 109 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_data_in[25]
port 110 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 la_data_in[26]
port 111 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_data_in[27]
port 112 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 la_data_in[28]
port 113 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_data_in[29]
port 114 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 la_data_in[2]
port 115 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 la_data_in[30]
port 116 nsew signal input
rlabel metal2 s 101310 0 101366 800 6 la_data_in[31]
port 117 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 la_data_in[32]
port 118 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 la_data_in[33]
port 119 nsew signal input
rlabel metal2 s 110418 0 110474 800 6 la_data_in[34]
port 120 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 la_data_in[35]
port 121 nsew signal input
rlabel metal2 s 116490 0 116546 800 6 la_data_in[36]
port 122 nsew signal input
rlabel metal2 s 119526 0 119582 800 6 la_data_in[37]
port 123 nsew signal input
rlabel metal2 s 122562 0 122618 800 6 la_data_in[38]
port 124 nsew signal input
rlabel metal2 s 125598 0 125654 800 6 la_data_in[39]
port 125 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 la_data_in[3]
port 126 nsew signal input
rlabel metal2 s 128634 0 128690 800 6 la_data_in[40]
port 127 nsew signal input
rlabel metal2 s 131670 0 131726 800 6 la_data_in[41]
port 128 nsew signal input
rlabel metal2 s 134706 0 134762 800 6 la_data_in[42]
port 129 nsew signal input
rlabel metal2 s 137742 0 137798 800 6 la_data_in[43]
port 130 nsew signal input
rlabel metal2 s 140778 0 140834 800 6 la_data_in[44]
port 131 nsew signal input
rlabel metal2 s 143814 0 143870 800 6 la_data_in[45]
port 132 nsew signal input
rlabel metal2 s 146850 0 146906 800 6 la_data_in[46]
port 133 nsew signal input
rlabel metal2 s 149886 0 149942 800 6 la_data_in[47]
port 134 nsew signal input
rlabel metal2 s 152922 0 152978 800 6 la_data_in[48]
port 135 nsew signal input
rlabel metal2 s 155958 0 156014 800 6 la_data_in[49]
port 136 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 la_data_in[4]
port 137 nsew signal input
rlabel metal2 s 158994 0 159050 800 6 la_data_in[50]
port 138 nsew signal input
rlabel metal2 s 162030 0 162086 800 6 la_data_in[51]
port 139 nsew signal input
rlabel metal2 s 165066 0 165122 800 6 la_data_in[52]
port 140 nsew signal input
rlabel metal2 s 168102 0 168158 800 6 la_data_in[53]
port 141 nsew signal input
rlabel metal2 s 171138 0 171194 800 6 la_data_in[54]
port 142 nsew signal input
rlabel metal2 s 174174 0 174230 800 6 la_data_in[55]
port 143 nsew signal input
rlabel metal2 s 177210 0 177266 800 6 la_data_in[56]
port 144 nsew signal input
rlabel metal2 s 180246 0 180302 800 6 la_data_in[57]
port 145 nsew signal input
rlabel metal2 s 183282 0 183338 800 6 la_data_in[58]
port 146 nsew signal input
rlabel metal2 s 186318 0 186374 800 6 la_data_in[59]
port 147 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 la_data_in[5]
port 148 nsew signal input
rlabel metal2 s 189354 0 189410 800 6 la_data_in[60]
port 149 nsew signal input
rlabel metal2 s 192390 0 192446 800 6 la_data_in[61]
port 150 nsew signal input
rlabel metal2 s 195426 0 195482 800 6 la_data_in[62]
port 151 nsew signal input
rlabel metal2 s 198462 0 198518 800 6 la_data_in[63]
port 152 nsew signal input
rlabel metal2 s 201498 0 201554 800 6 la_data_in[64]
port 153 nsew signal input
rlabel metal2 s 204534 0 204590 800 6 la_data_in[65]
port 154 nsew signal input
rlabel metal2 s 207570 0 207626 800 6 la_data_in[66]
port 155 nsew signal input
rlabel metal2 s 210606 0 210662 800 6 la_data_in[67]
port 156 nsew signal input
rlabel metal2 s 213642 0 213698 800 6 la_data_in[68]
port 157 nsew signal input
rlabel metal2 s 216678 0 216734 800 6 la_data_in[69]
port 158 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 la_data_in[6]
port 159 nsew signal input
rlabel metal2 s 219714 0 219770 800 6 la_data_in[70]
port 160 nsew signal input
rlabel metal2 s 222750 0 222806 800 6 la_data_in[71]
port 161 nsew signal input
rlabel metal2 s 225786 0 225842 800 6 la_data_in[72]
port 162 nsew signal input
rlabel metal2 s 228822 0 228878 800 6 la_data_in[73]
port 163 nsew signal input
rlabel metal2 s 231858 0 231914 800 6 la_data_in[74]
port 164 nsew signal input
rlabel metal2 s 234894 0 234950 800 6 la_data_in[75]
port 165 nsew signal input
rlabel metal2 s 237930 0 237986 800 6 la_data_in[76]
port 166 nsew signal input
rlabel metal2 s 240966 0 241022 800 6 la_data_in[77]
port 167 nsew signal input
rlabel metal2 s 244002 0 244058 800 6 la_data_in[78]
port 168 nsew signal input
rlabel metal2 s 247038 0 247094 800 6 la_data_in[79]
port 169 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 la_data_in[7]
port 170 nsew signal input
rlabel metal2 s 250074 0 250130 800 6 la_data_in[80]
port 171 nsew signal input
rlabel metal2 s 253110 0 253166 800 6 la_data_in[81]
port 172 nsew signal input
rlabel metal2 s 256146 0 256202 800 6 la_data_in[82]
port 173 nsew signal input
rlabel metal2 s 259182 0 259238 800 6 la_data_in[83]
port 174 nsew signal input
rlabel metal2 s 262218 0 262274 800 6 la_data_in[84]
port 175 nsew signal input
rlabel metal2 s 265254 0 265310 800 6 la_data_in[85]
port 176 nsew signal input
rlabel metal2 s 268290 0 268346 800 6 la_data_in[86]
port 177 nsew signal input
rlabel metal2 s 271326 0 271382 800 6 la_data_in[87]
port 178 nsew signal input
rlabel metal2 s 274362 0 274418 800 6 la_data_in[88]
port 179 nsew signal input
rlabel metal2 s 277398 0 277454 800 6 la_data_in[89]
port 180 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 la_data_in[8]
port 181 nsew signal input
rlabel metal2 s 280434 0 280490 800 6 la_data_in[90]
port 182 nsew signal input
rlabel metal2 s 283470 0 283526 800 6 la_data_in[91]
port 183 nsew signal input
rlabel metal2 s 286506 0 286562 800 6 la_data_in[92]
port 184 nsew signal input
rlabel metal2 s 289542 0 289598 800 6 la_data_in[93]
port 185 nsew signal input
rlabel metal2 s 292578 0 292634 800 6 la_data_in[94]
port 186 nsew signal input
rlabel metal2 s 295614 0 295670 800 6 la_data_in[95]
port 187 nsew signal input
rlabel metal2 s 298650 0 298706 800 6 la_data_in[96]
port 188 nsew signal input
rlabel metal2 s 301686 0 301742 800 6 la_data_in[97]
port 189 nsew signal input
rlabel metal2 s 304722 0 304778 800 6 la_data_in[98]
port 190 nsew signal input
rlabel metal2 s 307758 0 307814 800 6 la_data_in[99]
port 191 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 la_data_in[9]
port 192 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 la_data_out[0]
port 193 nsew signal output
rlabel metal2 s 311806 0 311862 800 6 la_data_out[100]
port 194 nsew signal output
rlabel metal2 s 314842 0 314898 800 6 la_data_out[101]
port 195 nsew signal output
rlabel metal2 s 317878 0 317934 800 6 la_data_out[102]
port 196 nsew signal output
rlabel metal2 s 320914 0 320970 800 6 la_data_out[103]
port 197 nsew signal output
rlabel metal2 s 323950 0 324006 800 6 la_data_out[104]
port 198 nsew signal output
rlabel metal2 s 326986 0 327042 800 6 la_data_out[105]
port 199 nsew signal output
rlabel metal2 s 330022 0 330078 800 6 la_data_out[106]
port 200 nsew signal output
rlabel metal2 s 333058 0 333114 800 6 la_data_out[107]
port 201 nsew signal output
rlabel metal2 s 336094 0 336150 800 6 la_data_out[108]
port 202 nsew signal output
rlabel metal2 s 339130 0 339186 800 6 la_data_out[109]
port 203 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 la_data_out[10]
port 204 nsew signal output
rlabel metal2 s 342166 0 342222 800 6 la_data_out[110]
port 205 nsew signal output
rlabel metal2 s 345202 0 345258 800 6 la_data_out[111]
port 206 nsew signal output
rlabel metal2 s 348238 0 348294 800 6 la_data_out[112]
port 207 nsew signal output
rlabel metal2 s 351274 0 351330 800 6 la_data_out[113]
port 208 nsew signal output
rlabel metal2 s 354310 0 354366 800 6 la_data_out[114]
port 209 nsew signal output
rlabel metal2 s 357346 0 357402 800 6 la_data_out[115]
port 210 nsew signal output
rlabel metal2 s 360382 0 360438 800 6 la_data_out[116]
port 211 nsew signal output
rlabel metal2 s 363418 0 363474 800 6 la_data_out[117]
port 212 nsew signal output
rlabel metal2 s 366454 0 366510 800 6 la_data_out[118]
port 213 nsew signal output
rlabel metal2 s 369490 0 369546 800 6 la_data_out[119]
port 214 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 la_data_out[11]
port 215 nsew signal output
rlabel metal2 s 372526 0 372582 800 6 la_data_out[120]
port 216 nsew signal output
rlabel metal2 s 375562 0 375618 800 6 la_data_out[121]
port 217 nsew signal output
rlabel metal2 s 378598 0 378654 800 6 la_data_out[122]
port 218 nsew signal output
rlabel metal2 s 381634 0 381690 800 6 la_data_out[123]
port 219 nsew signal output
rlabel metal2 s 384670 0 384726 800 6 la_data_out[124]
port 220 nsew signal output
rlabel metal2 s 387706 0 387762 800 6 la_data_out[125]
port 221 nsew signal output
rlabel metal2 s 390742 0 390798 800 6 la_data_out[126]
port 222 nsew signal output
rlabel metal2 s 393778 0 393834 800 6 la_data_out[127]
port 223 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 la_data_out[12]
port 224 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 la_data_out[13]
port 225 nsew signal output
rlabel metal2 s 50710 0 50766 800 6 la_data_out[14]
port 226 nsew signal output
rlabel metal2 s 53746 0 53802 800 6 la_data_out[15]
port 227 nsew signal output
rlabel metal2 s 56782 0 56838 800 6 la_data_out[16]
port 228 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 la_data_out[17]
port 229 nsew signal output
rlabel metal2 s 62854 0 62910 800 6 la_data_out[18]
port 230 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 la_data_out[19]
port 231 nsew signal output
rlabel metal2 s 11242 0 11298 800 6 la_data_out[1]
port 232 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 la_data_out[20]
port 233 nsew signal output
rlabel metal2 s 71962 0 72018 800 6 la_data_out[21]
port 234 nsew signal output
rlabel metal2 s 74998 0 75054 800 6 la_data_out[22]
port 235 nsew signal output
rlabel metal2 s 78034 0 78090 800 6 la_data_out[23]
port 236 nsew signal output
rlabel metal2 s 81070 0 81126 800 6 la_data_out[24]
port 237 nsew signal output
rlabel metal2 s 84106 0 84162 800 6 la_data_out[25]
port 238 nsew signal output
rlabel metal2 s 87142 0 87198 800 6 la_data_out[26]
port 239 nsew signal output
rlabel metal2 s 90178 0 90234 800 6 la_data_out[27]
port 240 nsew signal output
rlabel metal2 s 93214 0 93270 800 6 la_data_out[28]
port 241 nsew signal output
rlabel metal2 s 96250 0 96306 800 6 la_data_out[29]
port 242 nsew signal output
rlabel metal2 s 14278 0 14334 800 6 la_data_out[2]
port 243 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 la_data_out[30]
port 244 nsew signal output
rlabel metal2 s 102322 0 102378 800 6 la_data_out[31]
port 245 nsew signal output
rlabel metal2 s 105358 0 105414 800 6 la_data_out[32]
port 246 nsew signal output
rlabel metal2 s 108394 0 108450 800 6 la_data_out[33]
port 247 nsew signal output
rlabel metal2 s 111430 0 111486 800 6 la_data_out[34]
port 248 nsew signal output
rlabel metal2 s 114466 0 114522 800 6 la_data_out[35]
port 249 nsew signal output
rlabel metal2 s 117502 0 117558 800 6 la_data_out[36]
port 250 nsew signal output
rlabel metal2 s 120538 0 120594 800 6 la_data_out[37]
port 251 nsew signal output
rlabel metal2 s 123574 0 123630 800 6 la_data_out[38]
port 252 nsew signal output
rlabel metal2 s 126610 0 126666 800 6 la_data_out[39]
port 253 nsew signal output
rlabel metal2 s 17314 0 17370 800 6 la_data_out[3]
port 254 nsew signal output
rlabel metal2 s 129646 0 129702 800 6 la_data_out[40]
port 255 nsew signal output
rlabel metal2 s 132682 0 132738 800 6 la_data_out[41]
port 256 nsew signal output
rlabel metal2 s 135718 0 135774 800 6 la_data_out[42]
port 257 nsew signal output
rlabel metal2 s 138754 0 138810 800 6 la_data_out[43]
port 258 nsew signal output
rlabel metal2 s 141790 0 141846 800 6 la_data_out[44]
port 259 nsew signal output
rlabel metal2 s 144826 0 144882 800 6 la_data_out[45]
port 260 nsew signal output
rlabel metal2 s 147862 0 147918 800 6 la_data_out[46]
port 261 nsew signal output
rlabel metal2 s 150898 0 150954 800 6 la_data_out[47]
port 262 nsew signal output
rlabel metal2 s 153934 0 153990 800 6 la_data_out[48]
port 263 nsew signal output
rlabel metal2 s 156970 0 157026 800 6 la_data_out[49]
port 264 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 la_data_out[4]
port 265 nsew signal output
rlabel metal2 s 160006 0 160062 800 6 la_data_out[50]
port 266 nsew signal output
rlabel metal2 s 163042 0 163098 800 6 la_data_out[51]
port 267 nsew signal output
rlabel metal2 s 166078 0 166134 800 6 la_data_out[52]
port 268 nsew signal output
rlabel metal2 s 169114 0 169170 800 6 la_data_out[53]
port 269 nsew signal output
rlabel metal2 s 172150 0 172206 800 6 la_data_out[54]
port 270 nsew signal output
rlabel metal2 s 175186 0 175242 800 6 la_data_out[55]
port 271 nsew signal output
rlabel metal2 s 178222 0 178278 800 6 la_data_out[56]
port 272 nsew signal output
rlabel metal2 s 181258 0 181314 800 6 la_data_out[57]
port 273 nsew signal output
rlabel metal2 s 184294 0 184350 800 6 la_data_out[58]
port 274 nsew signal output
rlabel metal2 s 187330 0 187386 800 6 la_data_out[59]
port 275 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 la_data_out[5]
port 276 nsew signal output
rlabel metal2 s 190366 0 190422 800 6 la_data_out[60]
port 277 nsew signal output
rlabel metal2 s 193402 0 193458 800 6 la_data_out[61]
port 278 nsew signal output
rlabel metal2 s 196438 0 196494 800 6 la_data_out[62]
port 279 nsew signal output
rlabel metal2 s 199474 0 199530 800 6 la_data_out[63]
port 280 nsew signal output
rlabel metal2 s 202510 0 202566 800 6 la_data_out[64]
port 281 nsew signal output
rlabel metal2 s 205546 0 205602 800 6 la_data_out[65]
port 282 nsew signal output
rlabel metal2 s 208582 0 208638 800 6 la_data_out[66]
port 283 nsew signal output
rlabel metal2 s 211618 0 211674 800 6 la_data_out[67]
port 284 nsew signal output
rlabel metal2 s 214654 0 214710 800 6 la_data_out[68]
port 285 nsew signal output
rlabel metal2 s 217690 0 217746 800 6 la_data_out[69]
port 286 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 la_data_out[6]
port 287 nsew signal output
rlabel metal2 s 220726 0 220782 800 6 la_data_out[70]
port 288 nsew signal output
rlabel metal2 s 223762 0 223818 800 6 la_data_out[71]
port 289 nsew signal output
rlabel metal2 s 226798 0 226854 800 6 la_data_out[72]
port 290 nsew signal output
rlabel metal2 s 229834 0 229890 800 6 la_data_out[73]
port 291 nsew signal output
rlabel metal2 s 232870 0 232926 800 6 la_data_out[74]
port 292 nsew signal output
rlabel metal2 s 235906 0 235962 800 6 la_data_out[75]
port 293 nsew signal output
rlabel metal2 s 238942 0 238998 800 6 la_data_out[76]
port 294 nsew signal output
rlabel metal2 s 241978 0 242034 800 6 la_data_out[77]
port 295 nsew signal output
rlabel metal2 s 245014 0 245070 800 6 la_data_out[78]
port 296 nsew signal output
rlabel metal2 s 248050 0 248106 800 6 la_data_out[79]
port 297 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 la_data_out[7]
port 298 nsew signal output
rlabel metal2 s 251086 0 251142 800 6 la_data_out[80]
port 299 nsew signal output
rlabel metal2 s 254122 0 254178 800 6 la_data_out[81]
port 300 nsew signal output
rlabel metal2 s 257158 0 257214 800 6 la_data_out[82]
port 301 nsew signal output
rlabel metal2 s 260194 0 260250 800 6 la_data_out[83]
port 302 nsew signal output
rlabel metal2 s 263230 0 263286 800 6 la_data_out[84]
port 303 nsew signal output
rlabel metal2 s 266266 0 266322 800 6 la_data_out[85]
port 304 nsew signal output
rlabel metal2 s 269302 0 269358 800 6 la_data_out[86]
port 305 nsew signal output
rlabel metal2 s 272338 0 272394 800 6 la_data_out[87]
port 306 nsew signal output
rlabel metal2 s 275374 0 275430 800 6 la_data_out[88]
port 307 nsew signal output
rlabel metal2 s 278410 0 278466 800 6 la_data_out[89]
port 308 nsew signal output
rlabel metal2 s 32494 0 32550 800 6 la_data_out[8]
port 309 nsew signal output
rlabel metal2 s 281446 0 281502 800 6 la_data_out[90]
port 310 nsew signal output
rlabel metal2 s 284482 0 284538 800 6 la_data_out[91]
port 311 nsew signal output
rlabel metal2 s 287518 0 287574 800 6 la_data_out[92]
port 312 nsew signal output
rlabel metal2 s 290554 0 290610 800 6 la_data_out[93]
port 313 nsew signal output
rlabel metal2 s 293590 0 293646 800 6 la_data_out[94]
port 314 nsew signal output
rlabel metal2 s 296626 0 296682 800 6 la_data_out[95]
port 315 nsew signal output
rlabel metal2 s 299662 0 299718 800 6 la_data_out[96]
port 316 nsew signal output
rlabel metal2 s 302698 0 302754 800 6 la_data_out[97]
port 317 nsew signal output
rlabel metal2 s 305734 0 305790 800 6 la_data_out[98]
port 318 nsew signal output
rlabel metal2 s 308770 0 308826 800 6 la_data_out[99]
port 319 nsew signal output
rlabel metal2 s 35530 0 35586 800 6 la_data_out[9]
port 320 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 la_oenb[0]
port 321 nsew signal input
rlabel metal2 s 312818 0 312874 800 6 la_oenb[100]
port 322 nsew signal input
rlabel metal2 s 315854 0 315910 800 6 la_oenb[101]
port 323 nsew signal input
rlabel metal2 s 318890 0 318946 800 6 la_oenb[102]
port 324 nsew signal input
rlabel metal2 s 321926 0 321982 800 6 la_oenb[103]
port 325 nsew signal input
rlabel metal2 s 324962 0 325018 800 6 la_oenb[104]
port 326 nsew signal input
rlabel metal2 s 327998 0 328054 800 6 la_oenb[105]
port 327 nsew signal input
rlabel metal2 s 331034 0 331090 800 6 la_oenb[106]
port 328 nsew signal input
rlabel metal2 s 334070 0 334126 800 6 la_oenb[107]
port 329 nsew signal input
rlabel metal2 s 337106 0 337162 800 6 la_oenb[108]
port 330 nsew signal input
rlabel metal2 s 340142 0 340198 800 6 la_oenb[109]
port 331 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 la_oenb[10]
port 332 nsew signal input
rlabel metal2 s 343178 0 343234 800 6 la_oenb[110]
port 333 nsew signal input
rlabel metal2 s 346214 0 346270 800 6 la_oenb[111]
port 334 nsew signal input
rlabel metal2 s 349250 0 349306 800 6 la_oenb[112]
port 335 nsew signal input
rlabel metal2 s 352286 0 352342 800 6 la_oenb[113]
port 336 nsew signal input
rlabel metal2 s 355322 0 355378 800 6 la_oenb[114]
port 337 nsew signal input
rlabel metal2 s 358358 0 358414 800 6 la_oenb[115]
port 338 nsew signal input
rlabel metal2 s 361394 0 361450 800 6 la_oenb[116]
port 339 nsew signal input
rlabel metal2 s 364430 0 364486 800 6 la_oenb[117]
port 340 nsew signal input
rlabel metal2 s 367466 0 367522 800 6 la_oenb[118]
port 341 nsew signal input
rlabel metal2 s 370502 0 370558 800 6 la_oenb[119]
port 342 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 la_oenb[11]
port 343 nsew signal input
rlabel metal2 s 373538 0 373594 800 6 la_oenb[120]
port 344 nsew signal input
rlabel metal2 s 376574 0 376630 800 6 la_oenb[121]
port 345 nsew signal input
rlabel metal2 s 379610 0 379666 800 6 la_oenb[122]
port 346 nsew signal input
rlabel metal2 s 382646 0 382702 800 6 la_oenb[123]
port 347 nsew signal input
rlabel metal2 s 385682 0 385738 800 6 la_oenb[124]
port 348 nsew signal input
rlabel metal2 s 388718 0 388774 800 6 la_oenb[125]
port 349 nsew signal input
rlabel metal2 s 391754 0 391810 800 6 la_oenb[126]
port 350 nsew signal input
rlabel metal2 s 394790 0 394846 800 6 la_oenb[127]
port 351 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 la_oenb[12]
port 352 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 la_oenb[13]
port 353 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 la_oenb[14]
port 354 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 la_oenb[15]
port 355 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_oenb[16]
port 356 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 la_oenb[17]
port 357 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_oenb[18]
port 358 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 la_oenb[19]
port 359 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 la_oenb[1]
port 360 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 la_oenb[20]
port 361 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_oenb[21]
port 362 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_oenb[22]
port 363 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 la_oenb[23]
port 364 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 la_oenb[24]
port 365 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_oenb[25]
port 366 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 la_oenb[26]
port 367 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 la_oenb[27]
port 368 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_oenb[28]
port 369 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_oenb[29]
port 370 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 la_oenb[2]
port 371 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 la_oenb[30]
port 372 nsew signal input
rlabel metal2 s 103334 0 103390 800 6 la_oenb[31]
port 373 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 la_oenb[32]
port 374 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 la_oenb[33]
port 375 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 la_oenb[34]
port 376 nsew signal input
rlabel metal2 s 115478 0 115534 800 6 la_oenb[35]
port 377 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 la_oenb[36]
port 378 nsew signal input
rlabel metal2 s 121550 0 121606 800 6 la_oenb[37]
port 379 nsew signal input
rlabel metal2 s 124586 0 124642 800 6 la_oenb[38]
port 380 nsew signal input
rlabel metal2 s 127622 0 127678 800 6 la_oenb[39]
port 381 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 la_oenb[3]
port 382 nsew signal input
rlabel metal2 s 130658 0 130714 800 6 la_oenb[40]
port 383 nsew signal input
rlabel metal2 s 133694 0 133750 800 6 la_oenb[41]
port 384 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 la_oenb[42]
port 385 nsew signal input
rlabel metal2 s 139766 0 139822 800 6 la_oenb[43]
port 386 nsew signal input
rlabel metal2 s 142802 0 142858 800 6 la_oenb[44]
port 387 nsew signal input
rlabel metal2 s 145838 0 145894 800 6 la_oenb[45]
port 388 nsew signal input
rlabel metal2 s 148874 0 148930 800 6 la_oenb[46]
port 389 nsew signal input
rlabel metal2 s 151910 0 151966 800 6 la_oenb[47]
port 390 nsew signal input
rlabel metal2 s 154946 0 155002 800 6 la_oenb[48]
port 391 nsew signal input
rlabel metal2 s 157982 0 158038 800 6 la_oenb[49]
port 392 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 la_oenb[4]
port 393 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 la_oenb[50]
port 394 nsew signal input
rlabel metal2 s 164054 0 164110 800 6 la_oenb[51]
port 395 nsew signal input
rlabel metal2 s 167090 0 167146 800 6 la_oenb[52]
port 396 nsew signal input
rlabel metal2 s 170126 0 170182 800 6 la_oenb[53]
port 397 nsew signal input
rlabel metal2 s 173162 0 173218 800 6 la_oenb[54]
port 398 nsew signal input
rlabel metal2 s 176198 0 176254 800 6 la_oenb[55]
port 399 nsew signal input
rlabel metal2 s 179234 0 179290 800 6 la_oenb[56]
port 400 nsew signal input
rlabel metal2 s 182270 0 182326 800 6 la_oenb[57]
port 401 nsew signal input
rlabel metal2 s 185306 0 185362 800 6 la_oenb[58]
port 402 nsew signal input
rlabel metal2 s 188342 0 188398 800 6 la_oenb[59]
port 403 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 la_oenb[5]
port 404 nsew signal input
rlabel metal2 s 191378 0 191434 800 6 la_oenb[60]
port 405 nsew signal input
rlabel metal2 s 194414 0 194470 800 6 la_oenb[61]
port 406 nsew signal input
rlabel metal2 s 197450 0 197506 800 6 la_oenb[62]
port 407 nsew signal input
rlabel metal2 s 200486 0 200542 800 6 la_oenb[63]
port 408 nsew signal input
rlabel metal2 s 203522 0 203578 800 6 la_oenb[64]
port 409 nsew signal input
rlabel metal2 s 206558 0 206614 800 6 la_oenb[65]
port 410 nsew signal input
rlabel metal2 s 209594 0 209650 800 6 la_oenb[66]
port 411 nsew signal input
rlabel metal2 s 212630 0 212686 800 6 la_oenb[67]
port 412 nsew signal input
rlabel metal2 s 215666 0 215722 800 6 la_oenb[68]
port 413 nsew signal input
rlabel metal2 s 218702 0 218758 800 6 la_oenb[69]
port 414 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 la_oenb[6]
port 415 nsew signal input
rlabel metal2 s 221738 0 221794 800 6 la_oenb[70]
port 416 nsew signal input
rlabel metal2 s 224774 0 224830 800 6 la_oenb[71]
port 417 nsew signal input
rlabel metal2 s 227810 0 227866 800 6 la_oenb[72]
port 418 nsew signal input
rlabel metal2 s 230846 0 230902 800 6 la_oenb[73]
port 419 nsew signal input
rlabel metal2 s 233882 0 233938 800 6 la_oenb[74]
port 420 nsew signal input
rlabel metal2 s 236918 0 236974 800 6 la_oenb[75]
port 421 nsew signal input
rlabel metal2 s 239954 0 240010 800 6 la_oenb[76]
port 422 nsew signal input
rlabel metal2 s 242990 0 243046 800 6 la_oenb[77]
port 423 nsew signal input
rlabel metal2 s 246026 0 246082 800 6 la_oenb[78]
port 424 nsew signal input
rlabel metal2 s 249062 0 249118 800 6 la_oenb[79]
port 425 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 la_oenb[7]
port 426 nsew signal input
rlabel metal2 s 252098 0 252154 800 6 la_oenb[80]
port 427 nsew signal input
rlabel metal2 s 255134 0 255190 800 6 la_oenb[81]
port 428 nsew signal input
rlabel metal2 s 258170 0 258226 800 6 la_oenb[82]
port 429 nsew signal input
rlabel metal2 s 261206 0 261262 800 6 la_oenb[83]
port 430 nsew signal input
rlabel metal2 s 264242 0 264298 800 6 la_oenb[84]
port 431 nsew signal input
rlabel metal2 s 267278 0 267334 800 6 la_oenb[85]
port 432 nsew signal input
rlabel metal2 s 270314 0 270370 800 6 la_oenb[86]
port 433 nsew signal input
rlabel metal2 s 273350 0 273406 800 6 la_oenb[87]
port 434 nsew signal input
rlabel metal2 s 276386 0 276442 800 6 la_oenb[88]
port 435 nsew signal input
rlabel metal2 s 279422 0 279478 800 6 la_oenb[89]
port 436 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 la_oenb[8]
port 437 nsew signal input
rlabel metal2 s 282458 0 282514 800 6 la_oenb[90]
port 438 nsew signal input
rlabel metal2 s 285494 0 285550 800 6 la_oenb[91]
port 439 nsew signal input
rlabel metal2 s 288530 0 288586 800 6 la_oenb[92]
port 440 nsew signal input
rlabel metal2 s 291566 0 291622 800 6 la_oenb[93]
port 441 nsew signal input
rlabel metal2 s 294602 0 294658 800 6 la_oenb[94]
port 442 nsew signal input
rlabel metal2 s 297638 0 297694 800 6 la_oenb[95]
port 443 nsew signal input
rlabel metal2 s 300674 0 300730 800 6 la_oenb[96]
port 444 nsew signal input
rlabel metal2 s 303710 0 303766 800 6 la_oenb[97]
port 445 nsew signal input
rlabel metal2 s 306746 0 306802 800 6 la_oenb[98]
port 446 nsew signal input
rlabel metal2 s 309782 0 309838 800 6 la_oenb[99]
port 447 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_oenb[9]
port 448 nsew signal input
rlabel metal4 s 4208 2128 4528 497808 6 vccd1
port 449 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 497808 6 vccd1
port 449 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 497808 6 vccd1
port 449 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 497808 6 vccd1
port 449 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 497808 6 vccd1
port 449 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 497808 6 vccd1
port 449 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 497808 6 vccd1
port 449 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 497808 6 vccd1
port 449 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 497808 6 vccd1
port 449 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 497808 6 vccd1
port 449 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 497808 6 vccd1
port 449 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 497808 6 vccd1
port 449 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 497808 6 vccd1
port 449 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 497808 6 vssd1
port 450 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 497808 6 vssd1
port 450 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 497808 6 vssd1
port 450 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 497808 6 vssd1
port 450 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 497808 6 vssd1
port 450 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 497808 6 vssd1
port 450 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 497808 6 vssd1
port 450 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 497808 6 vssd1
port 450 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 497808 6 vssd1
port 450 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 497808 6 vssd1
port 450 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 497808 6 vssd1
port 450 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 497808 6 vssd1
port 450 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 497808 6 vssd1
port 450 nsew ground bidirectional
rlabel metal2 s 5170 0 5226 800 6 wb_clk_i
port 451 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wb_rst_i
port 452 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 400000 500000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 75029958
string GDS_FILE /home/nick/sdmay25-28/openlane/user_proj_datapath/runs/24_10_31_23_47/results/signoff/user_proj_datapath.magic.gds
string GDS_START 545438
<< end >>

